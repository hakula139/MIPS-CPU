`ifndef BPB_SVH
`define BPB_SVH

`timescale 1ns / 1ps

// number of entries
`define BPB_E 8
// index bits
`define BPB_T 10

`endif
