`ifndef CACHE_CONTROLLER_SVH
`define CACHE_CONTROLLER_SVH

`define STATE_WIDTH 2

`define INITIAL    2'b00
`define WRITE_BACK 2'b01
`define READ_MEM   2'b10
`define ONLY_WRITE 2'b11

`endif
