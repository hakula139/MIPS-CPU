`ifndef CACHE_CONTROLLER_VH
`define CACHE_CONTROLLER_VH

`define STATE_WIDTH 2

`define INITIAL    2'b00
`define WRITE_BACK 2'b01
`define READ_MEM   2'b10

`endif