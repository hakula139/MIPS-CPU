`ifndef REPLACE_CONTROLLER_SVH
`define REPLACE_CONTROLLER_SVH

`define MODE_WIDTH 3

`define LRU 0
`define RR  1
`define LFU 2

`define REPLACE_MODE `LRU

`endif
