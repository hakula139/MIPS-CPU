`ifndef REPLACE_CONTROLLER_SVH
`define REPLACE_CONTROLLER_SVH

`define LRU 0
`define RR  1

`define REPLACE_MODE `LRU

`endif
